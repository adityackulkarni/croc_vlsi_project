// This module is supposed to issue one write transaction via OBI to SRAM0.
// Will require internal FSM.

module obi_writer (
    ports
);
    
endmodule