// This module is supposed to issue 8 read transactions via OBI to SRAM0. 
// Will require internal FSM.

module obi_reader (

)

endmodule
