// Copyright 2024 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Authors:
// - Philippe Sauter <phsauter@iis.ee.ethz.ch>

module user_domain import user_pkg::*; import croc_pkg::*; #(
  parameter int unsigned GpioCount = 16
) (
  input  logic      clk_i,
  input  logic      ref_clk_i,
  input  logic      rst_ni,
  input  logic      testmode_i,
  
  input  sbr_obi_req_t user_sbr_obi_req_i, // User Sbr (rsp_o), Croc Mgr (req_i)
  output sbr_obi_rsp_t user_sbr_obi_rsp_o,

  output mgr_obi_req_t user_mgr_obi_req_o, // User Mgr (req_o), Croc Sbr (rsp_i)
  input  mgr_obi_rsp_t user_mgr_obi_rsp_i,

  input  logic [      GpioCount-1:0] gpio_in_sync_i, // synchronized GPIO inputs
  output logic [NumExternalIrqs-1:0] interrupts_o // interrupts to core
);

  assign interrupts_o = '0;  


  //////////////////////
  // User Manager MUX //
  /////////////////////

  // No manager so we don't need a obi_mux module and just terminate the request properly
  assign user_mgr_obi_req_o = '0;


  ////////////////////////////
  // User Subordinate DEMUX //
  ////////////////////////////

  // ----------------------------------------------------------------------------------------------
  // User Subordinate Buses
  // ----------------------------------------------------------------------------------------------
  
  // collection of signals from the demultiplexer
  sbr_obi_req_t [NumDemuxSbr-1:0] all_user_sbr_obi_req;
  sbr_obi_rsp_t [NumDemuxSbr-1:0] all_user_sbr_obi_rsp;

  // Error Subordinate Bus
  sbr_obi_req_t user_error_obi_req;
  sbr_obi_rsp_t user_error_obi_rsp;

  // Fanout into more readable signals
  assign user_error_obi_req              = all_user_sbr_obi_req[UserError];
  assign all_user_sbr_obi_rsp[UserError] = user_error_obi_rsp;

  
  // Change - 6:
  // MMIO control signals from/to tbd_accel
  logic start_reg;
  logic done_reg;
  logic match_reg;


  // Change - 4:

  // Accelerator subordinate (tbd_accel)
  sbr_obi_req_t user_tbd_obi_req;
  sbr_obi_rsp_t user_tbd_obi_rsp;

  assign user_tbd_obi_req              = all_user_sbr_obi_req[UserTbd];
  // UserTbd is defined in user_pkg.sv
  assign all_user_sbr_obi_rsp[UserTbd] = user_tbd_obi_rsp;



  //-----------------------------------------------------------------------------------------------
  // Demultiplex to User Subordinates according to address map
  //-----------------------------------------------------------------------------------------------

  logic [cf_math_pkg::idx_width(NumDemuxSbr)-1:0] user_idx;

  addr_decode #(
    .NoIndices ( NumDemuxSbr                    ),
    .NoRules   ( NumDemuxSbrRules               ),
    .addr_t    ( logic[SbrObiCfg.DataWidth-1:0] ),
    .rule_t    ( addr_map_rule_t                ),
    .Napot     ( 1'b0                           )
  ) i_addr_decode_periphs (
    .addr_i           ( user_sbr_obi_req_i.a.addr ),
    .addr_map_i       ( user_addr_map             ),
    .idx_o            ( user_idx                  ),
    .dec_valid_o      (),
    .dec_error_o      (),
    .en_default_idx_i ( 1'b1 ),
    .default_idx_i    ( '0   )
  );

  obi_demux #(
    .ObiCfg      ( SbrObiCfg     ),
    .obi_req_t   ( sbr_obi_req_t ),
    .obi_rsp_t   ( sbr_obi_rsp_t ),
    .NumMgrPorts ( NumDemuxSbr   ),
    .NumMaxTrans ( 2             )
  ) i_obi_demux (
    .clk_i,
    .rst_ni,

    .sbr_port_select_i ( user_idx             ),
    .sbr_port_req_i    ( user_sbr_obi_req_i   ),
    .sbr_port_rsp_o    ( user_sbr_obi_rsp_o   ),

    .mgr_ports_req_o   ( all_user_sbr_obi_req ),
    .mgr_ports_rsp_i   ( all_user_sbr_obi_rsp )
  );


//-------------------------------------------------------------------------------------------------
// User Subordinates
//-------------------------------------------------------------------------------------------------

  // Error Subordinate
  obi_err_sbr #(
    .ObiCfg      ( SbrObiCfg     ),
    .obi_req_t   ( sbr_obi_req_t ),
    .obi_rsp_t   ( sbr_obi_rsp_t ),
    .NumMaxTrans ( 1             ),
    .RspData     ( 32'hBADCAB1E  )
  ) i_user_err (
    .clk_i,
    .rst_ni,
    .testmode_i ( testmode_i      ),
    .obi_req_i  ( user_error_obi_req ),
    .obi_rsp_o  ( user_error_obi_rsp )
  );


  // Change - 7:

  // Simple module to map start/done/match to MMIO registers

  // Simple OBI MMIO register interface for tbd_accel
  obi_simple_mmio #(
    .ObiCfg     ( SbrObiCfg ),
    .DataWidth  ( 32        )
  ) i_tbd_accel_mmio (
    .clk_i,
    .rst_ni,
    .obi_req_i ( user_tbd_obi_req ),
    .obi_rsp_o ( user_tbd_obi_rsp ),

    // Register-mapped outputs to accelerator
    .start_o ( start_reg ),
    .done_i  ( done_reg  ),
    .match_i ( match_reg )
  );


  // Change - 5:
  // Instantiate tbd_accel:

  // Connecting it to the system-wide OBI bus
  // Giving it access to SRAM
  // Bringing it into the build

  tbd_accel #(
    .BASE_ADDR(32'h2000_0000)
  ) i_user_tbd_accel (
    .clk      ( clk_i        ),
    .rst_n    ( rst_ni       ),

    // SRAM interface
    .sram_addr   ( /* connect appropriately or leave unconnected for now */ ),
    .sram_req    ( /* connect appropriately or leave unconnected */ ),
    .sram_rdata  ( /* connect appropriately or leave unconnected */ ),
    .sram_rvalid ( /* connect appropriately or leave unconnected */ ),

    // MMIO interface via OBI bus (connect from demuxed req/rsp)
    .start ( user_tbd_obi_req.a.wdata[0] ), // Simple example: use wdata[0] as 'start'
    .done  ( /* optionally wire to a status register */ ),
    .match ( /* optionally wire to a status register */ )
  );


endmodule
